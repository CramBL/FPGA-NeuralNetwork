module Layer_4 #(parameter NN = 30, numWeight=784, dataWidth=16, layerNum=1, sigmoidSize=10, weightIntWidth=4, actType="relu")
    (
    input           clk,
    input           rst,
    input           weightValid,
    input           biasValid,
    input [31:0]    weightValue,
    input [31:0]    biasValue,
    input [31:0]    config_layer_num,
    input [31:0]    config_neuron_num,
    input           x_valid,
    input [dataWidth-1:0]    x_in,
    output [NN-1:0]     o_valid,
    output [NN*dataWidth-1:0]  x_out
    );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(0),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_0.mif"),.biasFile("b_4_0.mif"))n_0(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[0*dataWidth+:dataWidth]),
            .outvalid(o_valid[0])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(1),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_1.mif"),.biasFile("b_4_1.mif"))n_1(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[1*dataWidth+:dataWidth]),
            .outvalid(o_valid[1])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(2),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_2.mif"),.biasFile("b_4_2.mif"))n_2(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[2*dataWidth+:dataWidth]),
            .outvalid(o_valid[2])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(3),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_3.mif"),.biasFile("b_4_3.mif"))n_3(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[3*dataWidth+:dataWidth]),
            .outvalid(o_valid[3])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(4),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_4.mif"),.biasFile("b_4_4.mif"))n_4(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[4*dataWidth+:dataWidth]),
            .outvalid(o_valid[4])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(5),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_5.mif"),.biasFile("b_4_5.mif"))n_5(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[5*dataWidth+:dataWidth]),
            .outvalid(o_valid[5])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(6),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_6.mif"),.biasFile("b_4_6.mif"))n_6(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[6*dataWidth+:dataWidth]),
            .outvalid(o_valid[6])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(7),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_7.mif"),.biasFile("b_4_7.mif"))n_7(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[7*dataWidth+:dataWidth]),
            .outvalid(o_valid[7])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(8),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_8.mif"),.biasFile("b_4_8.mif"))n_8(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[8*dataWidth+:dataWidth]),
            .outvalid(o_valid[8])
            );
neuron #(.numWeight(numWeight),.layerNo(layerNum),.neuronNo(9),.dataWidth(dataWidth),.sigmoidSize(sigmoidSize),.weightIntWidth(weightIntWidth),.actType(actType),.weightFile("w_4_9.mif"),.biasFile("b_4_9.mif"))n_9(
            .clk(clk),
            .rst(rst),
            .myinput(x_in),
            .weightValid(weightValid),
            .biasValid(biasValid),
            .weightValue(weightValue),
            .biasValue(biasValue),
            .config_layer_num(config_layer_num),
            .config_neuron_num(config_neuron_num),
            .myinputValid(x_valid),
            .out(x_out[9*dataWidth+:dataWidth]),
            .outvalid(o_valid[9])
            );
endmodule